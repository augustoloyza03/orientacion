library verilog;
use verilog.vl_types.all;
entity ubicacion_vlg_vec_tst is
end ubicacion_vlg_vec_tst;
